module inst_mem(input [31:0]Address,output reg [31:0]inst);
reg [31:0] mem[0:1023];

initial begin
    
    mem[0]=32'b001000_00000_00001_0000000000101000;//addi R1 R0 40
    mem[1]=32'b001000_00000_00101_0000000000000000;//addi R5 R0 0
    mem[2]=32'b000100_00001_00000_0000000000000100;//beq R1 R0 END //LOOP
    mem[3]=32'b100011_00001_00100_0000001111100100;//lw  R4 996(R1)
    mem[4]=32'b000000_00101_00100_0010100000100000;//add R5 R4 R5
    mem[5]=32'b001000_00001_00001_1111111111111100;//addi R1 R1 -4
    mem[6]=32'b000011_00000_00000_0000000000000010;//J LOOP
    mem[7]=32'b101011_00000_00101_0000011111010000;//sw R5 2000(R0) //END
    
    //mem[0]=32'b000011_00000_00000_0000000000000100;//J LOOP
    //mem[1]=32'b001000_00001_00001_1111111111111100;//addi R1 R1 -4
    //mem[4]=32'b000000_11111_00000_0000000000001000;//Jr //LOOP

    //mem[0]=32'b000010_00000_00000_0000000000000011;//J LOOP

    //mem[3]=32'b001000_00001_00001_1111111111111100;//addi R1 R1 -4 //LOOP
    /*
    mem[0]=32'b001000_00000000010000000000101000;//addi R1 R0 40
    mem[1]=32'b001000_00001_00101_0000000000000000;//addi R5 R1 0
    mem[2]=32'b00000000101001000010100000100000;//add R5 R4 R5
    mem[3]=32'b100011_00001_00100_0000001111100100;//lw  R4 996(R1)
    mem[4]=32'b000000_00101_00100_0010100000100000;//add R5 R4 R5
    */
end

always @(Address) begin
    inst<=mem[Address[31:2]];
end
endmodule